netcdf parking_lot_photo_rates {

dimensions:
time = unlimited;

variables:
  double time(time);
  double O3_1(time);
  double O3_2(time);
  double O2_1(time);

  time:units = "hours";
  O3_1:units = "s-1";
  O3_2:units = "s-1";
  O2_1:units = "s-1";

}
